`ifndef AXIS_I2C_PKG
`define AXIS_I2C_PKG

package axis_i2c_pkg;

    parameter I2C_DATA_WIDTH  = 8;
    parameter I2C_ADDR_WIDTH  = 7;
    parameter AXIS_DATA_WIDTH = 16;
    parameter CNT_WIDTH       = $clog2(I2C_DATA_WIDTH);

endpackage

`endif
