interface axis_i2c_top_if;

    bit clk;
    bit arstn;

    logic i2c_sda;
    logic i2c_scl;

endinterface
